----------------------------------------------------------------------------------
-- TECHNICAL UNIVERSITY OF CRETE
-- NICK KYPARISSAS
-- MODULE: Toroidal Grid Lines Buffer, transmits a neighborhood column per clock cycle. 
-- PROJECT NAME: A Framework for the Real-Time Execution of Cellular Automata on Reconfigurable Logic
-- Diploma Thesis Project 2019
----------------------------------------------------------------------------------

-- VHDL 2008: FOR USING "PROCESS(ALL)"
	
-- GRID_LINES_TOROIDAL_BUFFER implements a toroidal grid consisting of 
-- GRID_X x GRID_Y cells. 
----------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY GRID_LINES_TOROIDAL_BUFFER IS
	GENERIC (
		CELL_SIZE : INTEGER := 4; 
		BURST_SIZE : INTEGER := 128;
		GRID_X : INTEGER := 1920;
		GRID_Y : INTEGER := 1080;
		NUMBER_OF_BURSTS_PER_LINE 	: INTEGER := 60; -- GRID_X * CELL_SIZE / BURST_SIZE;
		NEIGHBORHOOD_SIZE  	: INTEGER := 29;
		SPEED : INTEGER := 120); 
	PORT (
		CLK_200 : IN STD_LOGIC; -- SYSTEM CLOCK
		UI_CLK : IN STD_LOGIC; -- SYSTEM CLOCK
		RST_UI_CLK : IN STD_LOGIC; -- HIGH ACTIVE SYNCHRONOUS RESET
		RST_200	: IN STD_LOGIC;
		-- SIGNALS NEEDED FOR THE TOROIDAL GRID: 
		-- THE BUFFER NO LONGER WAITS FOR THE GRAPHICS FEEDER TO FEED IT!
		WRITE_BACK_COLUMN : IN INTEGER RANGE 0 TO NUMBER_OF_BURSTS_PER_LINE-1;
		WRITE_BACK_ROW : IN INTEGER RANGE 0 TO GRID_Y-1;
		INIT_COLUMN : IN INTEGER RANGE 0 TO NUMBER_OF_BURSTS_PER_LINE-1;
		INIT_ROW : IN INTEGER RANGE 0 TO GRID_Y-1;
		INIT_COMPLETE : IN STD_LOGIC; 
		SIM_ENDED : IN STD_LOGIC;
		SPEED_COUNTER : IN INTEGER RANGE 0 TO SPEED := 0;
		SPEED_SETTING : IN INTEGER RANGE 0 TO SPEED; -- GRAPHICS RUN AT 60 FPS. SPEED = 60: NEW GENERATION EVERY 1 SEC. SPEED = 0: FULL SPEED, NEW GENERATION EVERY NEW FRAME.
		--
		MEM_WRITE_DATA : IN STD_LOGIC_VECTOR(BURST_SIZE-1 DOWNTO 0);
		--APP_WDF_RDY : IN STD_LOGIC;
		APP_WDF_WREN : IN STD_LOGIC;
		-------------------
		WRITE_EN : IN STD_LOGIC;
		DATA_IN : IN STD_LOGIC_VECTOR(BURST_SIZE-1 DOWNTO 0);
		MEMORY_ACCESS_GRANTED : IN STD_LOGIC;
		DATA_OUT : OUT STD_LOGIC_VECTOR((NEIGHBORHOOD_SIZE*CELL_SIZE)-1 DOWNTO 0);
		DATA_OUT_VALID 	: OUT STD_LOGIC -- WHEN DATA_OUT_VALID = 1, THE ARRAY IS BEING DRAINED, ONE DATA_OUT COLUMN PER CLK CYCLE
		); 
END GRID_LINES_TOROIDAL_BUFFER;

ARCHITECTURE BEHAVIORAL OF GRID_LINES_TOROIDAL_BUFFER IS
	
	SIGNAL WRITE_ADDRESS_COUNTER : INTEGER RANGE 0 TO NUMBER_OF_BURSTS_PER_LINE-1 := 0;
	SIGNAL READ_ADDRESS_COUNTER : INTEGER RANGE 0 TO GRID_X-1 := GRID_X-((NEIGHBORHOOD_SIZE-1)/2);
	
	TYPE CRAPPY_SIGNAL IS ARRAY (NEIGHBORHOOD_SIZE+NEIGHBORHOOD_SIZE-1 DOWNTO 0) OF STD_LOGIC_VECTOR(0 DOWNTO 0); 
	SIGNAL WRITE_ENABLE : CRAPPY_SIGNAL := (OTHERS => (OTHERS => '0'));
	
	TYPE LINE_BUF_WRITE_SIG_TYPE IS ARRAY (NEIGHBORHOOD_SIZE+NEIGHBORHOOD_SIZE-1 DOWNTO 0) OF STD_LOGIC_VECTOR(6 DOWNTO 0);
	SIGNAL LINE_BUFFER_WR_ADDRESS, WRITE_ADDRESS : LINE_BUF_WRITE_SIG_TYPE;
	SIGNAL READ_ADDRESS : STD_LOGIC_VECTOR(10 DOWNTO 0);
	
	TYPE LINE_BUF_DATA_TYPE IS ARRAY (NEIGHBORHOOD_SIZE+NEIGHBORHOOD_SIZE-1 DOWNTO 0) OF STD_LOGIC_VECTOR(BURST_SIZE-1 DOWNTO 0);
	SIGNAL LINE_BUFFER_DATA_IN : LINE_BUF_DATA_TYPE;
	
	TYPE INTEGER_SYNCHRONIZER_1 IS ARRAY (1 DOWNTO 0) OF INTEGER RANGE 0 TO GRID_Y;
	SIGNAL TOTAL_NUM_OF_FILLED_LINES : INTEGER_SYNCHRONIZER_1;
	
	SIGNAL DATA_OUT_VALID_SIGNAL : STD_LOGIC_VECTOR(NEIGHBORHOOD_SIZE-1 DOWNTO 0) := (OTHERS => '0');
	
	TYPE INTEGER_SYNCHRONIZER_2 IS ARRAY (1 DOWNTO 0) OF INTEGER RANGE 0 TO NEIGHBORHOOD_SIZE;
	SIGNAL LINE_BEING_FILLED : INTEGER_SYNCHRONIZER_2;
	
	TYPE STD_LOGIC_ARRAY IS ARRAY (NEIGHBORHOOD_SIZE-1 DOWNTO 0, NEIGHBORHOOD_SIZE+NEIGHBORHOOD_SIZE-1 DOWNTO 0) OF STD_LOGIC_VECTOR(CELL_SIZE-1 DOWNTO 0);
	SIGNAL LINE_DATA : STD_LOGIC_ARRAY := (OTHERS => (OTHERS => (OTHERS => '0'))); 
	
	TYPE INTEGER_ARRAY IS ARRAY (NEIGHBORHOOD_SIZE-1 DOWNTO 0, NEIGHBORHOOD_SIZE-1 DOWNTO 0) OF INTEGER RANGE 0 TO NEIGHBORHOOD_SIZE+NEIGHBORHOOD_SIZE-1;
	SIGNAL LINES_BEING_DRAINED : INTEGER_ARRAY;
	SIGNAL LAST_LINE_BEING_DRAINED : INTEGER RANGE 0 TO NEIGHBORHOOD_SIZE;
	
	SIGNAL GRID_LINE_TO_BE_DRAINED : INTEGER RANGE 0 TO GRID_Y := 0; --((NEIGHBORHOOD_SIZE-1)/2);
	
	SIGNAL SYNC_CONTROL : STD_LOGIC := '0';
	
	TYPE STATE IS (RESET, WAIT_FOR_BUFFER_FILL, PRELOAD_NEIGHBORHOOD, BUFFER_DRAIN, WRAP_AROUND_NEIGHBORHOOD);
	SIGNAL FSM_STATE : STATE;	
	
	COMPONENT LINE_BUFFER_4b 
	PORT (
		clka : IN STD_LOGIC;
		wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
		addra : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		dina : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		clkb : IN STD_LOGIC;
		addrb : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		doutb : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
	END COMPONENT;
	
	COMPONENT LINE_BUFFER_8B 
	PORT (
		clka : IN STD_LOGIC;
		wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
		addra : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
		dina : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
		clkb : IN STD_LOGIC;
		addrb : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
		doutb : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
	END COMPONENT;
	-----------------------------------------------------
	constant BOUNDARY_CONDITION_01 : INTEGER := NEIGHBORHOOD_SIZE+((NEIGHBORHOOD_SIZE-1)/2)+1-(GRID_Y-1-(((NEIGHBORHOOD_SIZE-1)/2)-1)); 
	constant BOUNDARY_CONDITION_02 : INTEGER := GRID_Y-1-(((NEIGHBORHOOD_SIZE-1)/2)-1); 
	constant BOUNDARY_CONDITION_03 : INTEGER := GRID_Y-1;
	-----------------------------------------------------
	
BEGIN
		
	GENERATE_LINE_BUFFERS: for I in 0 to NEIGHBORHOOD_SIZE+NEIGHBORHOOD_SIZE-1 generate 
	-- 0 to NEIGHBORHOOD_SIZE-1 LINES + ONE FOR BUFFERING + NEIGHBORHOOD_SIZE-1 POLOIDAL BUFFERS
	-- 0 to NEIGHBORHOOD_SIZE for the common lines buffer
	-- NEIGHBORHOOD_SIZE+1 to NEIGHBORHOOD_SIZE+((NEIGHBORHOOD_SIZE-1)/2) for lines 0-2 (in 7x7)
	-- NEIGHBORHOOD_SIZE+((NEIGHBORHOOD_SIZE-1)/2)+1 to NEIGHBORHOOD_SIZE+NEIGHBORHOOD_SIZE-1 for lines 1077-1079 (in 7x7)
		LINE_BUFFER:	IF (CELL_SIZE = 4) GENERATE
			LINE_BUFFER_8: LINE_BUFFER_4b 
			PORT MAP(
				clka => UI_CLK,
				wea => WRITE_ENABLE(I),
				addra => LINE_BUFFER_WR_ADDRESS(I)(5 DOWNTO 0),
				dina => LINE_BUFFER_DATA_IN(I),
				clkb => CLK_200,
				addrb => READ_ADDRESS,
				doutb => LINE_DATA(0, I)
			); 
  		ELSIF (CELL_SIZE = 8) GENERATE
			LINE_BUFFER_8: LINE_BUFFER_8b 
			PORT MAP(
				clka => UI_CLK,
				wea => WRITE_ENABLE(I),
				addra => LINE_BUFFER_WR_ADDRESS(I),
				dina => LINE_BUFFER_DATA_IN(I),
				clkb => CLK_200,
				addrb => READ_ADDRESS,
				doutb => LINE_DATA(0, I)
			);
		END GENERATE LINE_BUFFER;
	end generate GENERATE_LINE_BUFFERS;
	
	SYNCHRONIZER: ENTITY WORK.SYNCHRONIZER
	GENERIC MAP (
		GRID_Y => GRID_Y,
		NEIGHBORHOOD_SIZE => NEIGHBORHOOD_SIZE
	) 
	PORT MAP (
		CLK_RX => CLK_200,
		RST => RST_200,
		--
		CONTROL => SYNC_CONTROL,
		DATA_IN_1 => TOTAL_NUM_OF_FILLED_LINES(0),
		DATA_OUT_1 => TOTAL_NUM_OF_FILLED_LINES(1),
		-- SYNCHRONIZING COMMUNICATING FSM SIGNALS:
		DATA_IN_2 => LINE_BEING_FILLED(0),
		DATA_OUT_2 => LINE_BEING_FILLED(1)
	);
	
	SET_BUFFER_SIGNALS: PROCESS(ALL) -- "PROCESS(ALL)" IS VHDL 2008!
	BEGIN
		for I in 0 to NEIGHBORHOOD_SIZE+NEIGHBORHOOD_SIZE-1 LOOP
			-- POLOIDAL_WRITE_ADDRESS <= STD_LOGIC_VECTOR(TO_UNSIGNED(WRITE_BACK_COLUMN, POLOIDAL_WRITE_ADDRESS'LENGTH)) WHEN INIT_COMPLETE = '1' ELSE STD_LOGIC_VECTOR(TO_UNSIGNED(INIT_COLUMN, POLOIDAL_WRITE_ADDRESS'LENGTH));
			-- WRITE_ADDRESS <= STD_LOGIC_VECTOR(TO_UNSIGNED(WRITE_ADDRESS_COUNTER, WRITE_ADDRESS'LENGTH));
			IF I >= NEIGHBORHOOD_SIZE+((NEIGHBORHOOD_SIZE-1)/2)+1 AND I <= NEIGHBORHOOD_SIZE+NEIGHBORHOOD_SIZE-1 THEN
				IF INIT_COMPLETE = '1' THEN 
					LINE_BUFFER_WR_ADDRESS(I) <= STD_LOGIC_VECTOR(TO_UNSIGNED(WRITE_BACK_COLUMN, LINE_BUFFER_WR_ADDRESS(I)'LENGTH));
				ELSE 
					LINE_BUFFER_WR_ADDRESS(I) <= STD_LOGIC_VECTOR(TO_UNSIGNED(INIT_COLUMN, LINE_BUFFER_WR_ADDRESS(I)'LENGTH));
				END IF;
				LINE_BUFFER_DATA_IN(I) <= MEM_WRITE_DATA;
			ELSE
				LINE_BUFFER_WR_ADDRESS(I) <= STD_LOGIC_VECTOR(TO_UNSIGNED(WRITE_ADDRESS_COUNTER, LINE_BUFFER_WR_ADDRESS(I)'LENGTH));
				LINE_BUFFER_DATA_IN(I) <= DATA_IN;
			END IF;
			
			-- SETTING WRITE_ENABLE
			IF I >= 0 AND I <= NEIGHBORHOOD_SIZE THEN
				IF I = LINE_BEING_FILLED(0) THEN
					WRITE_ENABLE(I)(0) <= WRITE_EN;
				ELSE
					WRITE_ENABLE(I)(0) <= '0';
				END IF;
			ELSIF I >= NEIGHBORHOOD_SIZE+1 AND I <= NEIGHBORHOOD_SIZE+((NEIGHBORHOOD_SIZE-1)/2) THEN
				-- THE FIRST LINES OF THE FRAME NEEDED FOR ITS CLOSURE COME FROM THE GRAPHICS FEEDER.
				-- HENCE, STRAIGHT FROM THE MEMORY. THE MEMORY CANT LET US KNOW WHICH LINE IT'S SENDING.
				-- THE LINE THAT'S COMING IS IDENTIFIED BY TOTAL_NUM_OF_FILLED_LINES. 
				IF I = LINE_BEING_FILLED(0) + NEIGHBORHOOD_SIZE + 1 AND TOTAL_NUM_OF_FILLED_LINES(0) < NEIGHBORHOOD_SIZE THEN
					WRITE_ENABLE(I)(0) <= WRITE_EN;
				ELSE
					WRITE_ENABLE(I)(0) <= '0';
				END IF;
			ELSE -- NEIGHBORHOOD_SIZE+((NEIGHBORHOOD_SIZE-1)/2)+1 to NEIGHBORHOOD_SIZE+NEIGHBORHOOD_SIZE-1 
				-- INIT AND WRITE-BACK LOAD THE BUFFER WITHT HE LAST LINES OF THE NEXT FRAME
				IF INIT_COMPLETE = '0' THEN
					-- IF LINE AT THE END OF THE FRAME WITHIN BOUNDARY CONDITIONS, ASSIGN IT TO THE RIGHT POLOIDAL BUFFER
					IF I = BOUNDARY_CONDITION_01+INIT_ROW AND INIT_ROW >= BOUNDARY_CONDITION_02 AND INIT_ROW <= BOUNDARY_CONDITION_03 THEN
						WRITE_ENABLE(I)(0) <= APP_WDF_WREN;
					ELSE
						WRITE_ENABLE(I) <= "0";
					END IF; 
				ELSE
					-- IF LINE AT THE END OF THE FRAME WITHIN BOUNDARY CONDITIONS, ASSIGN IT TO THE RIGHT POLOIDAL BUFFER
				IF I = BOUNDARY_CONDITION_01+WRITE_BACK_ROW AND WRITE_BACK_ROW >= BOUNDARY_CONDITION_02 AND WRITE_BACK_ROW <= BOUNDARY_CONDITION_03 AND SIM_ENDED = '0' AND SPEED_COUNTER >= SPEED_SETTING THEN 
						WRITE_ENABLE(I)(0) <= APP_WDF_WREN;
					ELSE
						WRITE_ENABLE(I) <= "0";
					END IF;	 
				END IF;
			END IF;
			
		END LOOP;
	END PROCESS;
	
	READ_ADDRESS <= STD_LOGIC_VECTOR(TO_UNSIGNED(READ_ADDRESS_COUNTER, READ_ADDRESS'LENGTH));
	

	
	WRITE: PROCESS
	BEGIN
		
		WAIT UNTIL RISING_EDGE(UI_CLK);		
		
		IF RST_UI_CLK = '1' THEN
			WRITE_ADDRESS_COUNTER <= 0;
			LINE_BEING_FILLED(0) <= 0;
			TOTAL_NUM_OF_FILLED_LINES(0) <= 0;
			SYNC_CONTROL <= '0';
		ELSE
			IF WRITE_EN = '1' AND MEMORY_ACCESS_GRANTED = '1' THEN
				IF WRITE_ADDRESS_COUNTER = NUMBER_OF_BURSTS_PER_LINE-1 THEN
					WRITE_ADDRESS_COUNTER <= 0;
					IF LINE_BEING_FILLED(0) = NEIGHBORHOOD_SIZE THEN 
					-- SOME SYNTHESIZERS WOULD CALCULATE THE OVERFLOW, BUT WE CHOOSE TO BE EXPLICIT
						LINE_BEING_FILLED(0) <= 0;
					ELSE
						LINE_BEING_FILLED(0) <= LINE_BEING_FILLED(0) + 1;
					END IF;
					-- NOTIFYING THE READER THERE IS A NEW LINE_BEING_FILLED VALUE
					TOTAL_NUM_OF_FILLED_LINES(0) <= TOTAL_NUM_OF_FILLED_LINES(0) + 1;
					SYNC_CONTROL <= '1';
				ELSE
					WRITE_ADDRESS_COUNTER <= WRITE_ADDRESS_COUNTER + 1;
					SYNC_CONTROL <= '0';
				END IF;
			ELSIF MEMORY_ACCESS_GRANTED = '0' AND TOTAL_NUM_OF_FILLED_LINES(0) = GRID_Y THEN
				-- NO ISSUE WITH COMMUNICATING WITH THE READING PROCESS:
				-- LINE_BEING_FILLED(0) <= 0; AFTER THAT PROCESS HAS STARTED DRAINING THE BUFFER
				TOTAL_NUM_OF_FILLED_LINES(0) <= 0;
				LINE_BEING_FILLED(0) <= 0;
				SYNC_CONTROL <= '1';
			ELSE 
				WRITE_ADDRESS_COUNTER <= WRITE_ADDRESS_COUNTER;
				TOTAL_NUM_OF_FILLED_LINES(0) <= TOTAL_NUM_OF_FILLED_LINES(0);
				LINE_BEING_FILLED(0) <= LINE_BEING_FILLED(0);
				SYNC_CONTROL <= '0';
			END IF;
		END IF;
	
	END PROCESS WRITE;

	
	READ: PROCESS
	BEGIN
		
		WAIT UNTIL RISING_EDGE(CLK_200);
		
		IF RST_200 = '1' THEN
			FSM_STATE <= RESET;
		ELSE
			CASE FSM_STATE IS 
			WHEN RESET =>
				FOR I IN 0 TO NEIGHBORHOOD_SIZE-1 LOOP
					IF I < ((NEIGHBORHOOD_SIZE-1)/2) THEN
						LINES_BEING_DRAINED(0, I) <= NEIGHBORHOOD_SIZE+((NEIGHBORHOOD_SIZE-1)/2)+1+I;
					ELSE
						LINES_BEING_DRAINED(0, I) <= I-((NEIGHBORHOOD_SIZE-1)/2); -- line 0 contains grid line (n-1) and so on 
						LAST_LINE_BEING_DRAINED <= I-((NEIGHBORHOOD_SIZE-1)/2); 
					END IF;
				END LOOP;
				GRID_LINE_TO_BE_DRAINED <= 0;
				READ_ADDRESS_COUNTER <= GRID_X-((NEIGHBORHOOD_SIZE-1)/2); -- RESET READ ADDRESS COUNTER
				DATA_OUT_VALID <= '0';
				DATA_OUT_VALID_SIGNAL <= (OTHERS => '0');
				FSM_STATE <= WAIT_FOR_BUFFER_FILL;
			WHEN WAIT_FOR_BUFFER_FILL => 
				IF (TOTAL_NUM_OF_FILLED_LINES(1) >= ((NEIGHBORHOOD_SIZE-1)/2)+1 AND LAST_LINE_BEING_DRAINED /= LINE_BEING_FILLED(1)) OR (GRID_LINE_TO_BE_DRAINED > GRID_Y-1-(NEIGHBORHOOD_SIZE/2) AND GRID_LINE_TO_BE_DRAINED < GRID_Y )  THEN  
					-- [ ((NEIGHBORHOOD_SIZE-1)/2)+1 ] + ((NEIGHBORHOOD_SIZE-1)/2) FROM THE POLOIDAL BUFFERS = NEIGHBORHOOD_SIZE
					-- IF THERE ARE ENOUGH LINES IN THE BUFFER 
					-- AND THE LINE WE ARE ABOUT TO DRAIN IS NOT THE ONE THAT'S BEING FILLED
					-- AND A NEW FRAME HAS BEEN LOADED
					-- OR IF WE ARE ABOUT TO WRAP AROUND POLOIDALLY THE GRID

					FSM_STATE <= PRELOAD_NEIGHBORHOOD;
				ELSE
					FSM_STATE <= FSM_STATE;  
				END IF;
				
				-- WE'RE APPROACHING THE END OF THE FRAME
				IF GRID_LINE_TO_BE_DRAINED = GRID_Y-1-(NEIGHBORHOOD_SIZE/2)+1 THEN
					LINES_BEING_DRAINED(0, NEIGHBORHOOD_SIZE-1) <= NEIGHBORHOOD_SIZE + 1;
				END IF;
				
				-- NEW FRAME: RESETTING WHICH LINES TO DRAIN
				-- IF TOTAL_NUM_OF_FILLED_LINES(1) = 0 THEN
				IF GRID_LINE_TO_BE_DRAINED = GRID_Y THEN
					FOR I IN 0 TO NEIGHBORHOOD_SIZE-1 LOOP
						IF I < ((NEIGHBORHOOD_SIZE-1)/2) THEN
							LINES_BEING_DRAINED(0, I) <= NEIGHBORHOOD_SIZE+((NEIGHBORHOOD_SIZE-1)/2)+1+I;
						ELSE
							LINES_BEING_DRAINED(0, I) <= I-((NEIGHBORHOOD_SIZE-1)/2); 
							LAST_LINE_BEING_DRAINED <= I-((NEIGHBORHOOD_SIZE-1)/2); 
						END IF;
					END LOOP; 
					GRID_LINE_TO_BE_DRAINED <= 0;
				END IF;
				
				DATA_OUT_VALID_SIGNAL(0) <= '0';
			
			WHEN PRELOAD_NEIGHBORHOOD =>
				
				IF READ_ADDRESS_COUNTER = GRID_X-1 THEN
					READ_ADDRESS_COUNTER <= 0;
				ELSE
					READ_ADDRESS_COUNTER <= READ_ADDRESS_COUNTER + 1;
				END IF;
				
				IF READ_ADDRESS_COUNTER = 0 THEN
					DATA_OUT_VALID_SIGNAL(0) <= '1';
					FSM_STATE <= BUFFER_DRAIN;
				ELSE
					FSM_STATE <= FSM_STATE;
				END IF;

			WHEN BUFFER_DRAIN => 
				 
				IF READ_ADDRESS_COUNTER = GRID_X-1 THEN
					READ_ADDRESS_COUNTER <= 0; 
					FSM_STATE <= WRAP_AROUND_NEIGHBORHOOD;  

				ELSE
					READ_ADDRESS_COUNTER <= READ_ADDRESS_COUNTER + 1;
					FSM_STATE <= FSM_STATE;
				END IF;
			
			WHEN WRAP_AROUND_NEIGHBORHOOD =>
				
				IF READ_ADDRESS_COUNTER = (NEIGHBORHOOD_SIZE-1)/2 THEN
					READ_ADDRESS_COUNTER <= GRID_X-((NEIGHBORHOOD_SIZE-1)/2); -- RESET READ ADDRESS COUNTER
					FOR I IN 0 TO NEIGHBORHOOD_SIZE-1 LOOP
						-- MOST SYNTHESIZERS WOULD CALCULATE THE OVERFLOW, BUT WE CHOOSE TO BE EXPLICIT
						IF LINES_BEING_DRAINED(0, I) = NEIGHBORHOOD_SIZE THEN
							LINES_BEING_DRAINED(0, I) <= 0;
						ELSE
							LINES_BEING_DRAINED(0, I) <= LINES_BEING_DRAINED(0, I) + 1;
						END IF; 
						IF LAST_LINE_BEING_DRAINED = NEIGHBORHOOD_SIZE THEN
							LAST_LINE_BEING_DRAINED <= 0;
						ELSE
							LAST_LINE_BEING_DRAINED <= LAST_LINE_BEING_DRAINED + 1;
						END IF; 
						-- GRADUALLY REPLACING THE LINES WINDOW WITH THE POLOIDAL BUFFER LINES 
						IF LINES_BEING_DRAINED(0, I) = NEIGHBORHOOD_SIZE + 1 AND I > 0 THEN
						-- IF WE'VE FOUND THE POLOIDAL WRAP-AROUND BUFFER (WHICH WILL BE NEIGHBORHOOD_SIZE + 2 AFTER THIS CYCLE), 
						-- THE PREVIOUS LINE OF THE WINDOW SHOULD BE REPLACED TO SLIDE DOWN
							LINES_BEING_DRAINED(0, I-1) <= LINES_BEING_DRAINED(0, I);
						END IF;
						-- SLIDING DOWN THE START OF THE FRAME
						IF LINES_BEING_DRAINED(0, I) = NEIGHBORHOOD_SIZE+(NEIGHBORHOOD_SIZE-1) AND I < NEIGHBORHOOD_SIZE-2 THEN
							LINES_BEING_DRAINED(0, I) <= LINES_BEING_DRAINED(0, I+1);
						END IF;
					END LOOP;
					
					GRID_LINE_TO_BE_DRAINED <= GRID_LINE_TO_BE_DRAINED + 1;
					
					FSM_STATE <= WAIT_FOR_BUFFER_FILL;
				ELSE
					READ_ADDRESS_COUNTER <= READ_ADDRESS_COUNTER + 1;
					FSM_STATE <= FSM_STATE;
				END IF;
				DATA_OUT_VALID_SIGNAL(0) <= '0';
				
			END CASE;
		END IF;
		
		-- PIPELINING REGISTERS FOR THE OUTPUTS
		-- AS THE SIZE OF NEIGHBORHOOD RISES, THE NUMBER OF BRAM MODULES RISES AS WELL
		-- ROUTING NEEDS MORE SLACK
		DATA_OUT_VALID <= DATA_OUT_VALID_SIGNAL(NEIGHBORHOOD_SIZE-1);
		FOR J IN NEIGHBORHOOD_SIZE-1 DOWNTO 1 LOOP	
			DATA_OUT_VALID_SIGNAL(J) <= DATA_OUT_VALID_SIGNAL(J-1);
		END LOOP;
		-- THE LINES BEING DRAINED CHANGE OVER TIME: (0, LINES_BEING_DRAINED(I))
		
		FOR I IN 0 TO NEIGHBORHOOD_SIZE-1 LOOP	
			DATA_OUT(((I+1)*CELL_SIZE)-1 DOWNTO (I*CELL_SIZE)) <= LINE_DATA(NEIGHBORHOOD_SIZE-1,  LINES_BEING_DRAINED(NEIGHBORHOOD_SIZE-1, I)); 
		END LOOP;
		
		L_1: FOR I IN 0 TO NEIGHBORHOOD_SIZE+NEIGHBORHOOD_SIZE-1 LOOP
			L_2: FOR J IN NEIGHBORHOOD_SIZE-1 DOWNTO 1 LOOP	
				LINE_DATA(J, I) <= LINE_DATA(J-1, I);
			END LOOP L_2;
		END LOOP L_1;
		
		L_3: FOR I IN 0 TO NEIGHBORHOOD_SIZE-1 LOOP
			L_4: FOR J IN NEIGHBORHOOD_SIZE-1 DOWNTO 1 LOOP	
				LINES_BEING_DRAINED(J, I) <= LINES_BEING_DRAINED(J-1, I);
			END LOOP L_4;
		END LOOP L_3;

	END PROCESS READ;
	
END BEHAVIORAL;