----------------------------------------------------------------------------------
-- TECHNICAL UNIVERSITY OF CRETE
-- NICK KYPARISSAS
-- MODULE: WRITE-BACK
-- PROJECT NAME: A Framework for the Real-Time Execution of Cellular Automata on Reconfigurable Logic
-- Diploma Thesis Project 2019
----------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY WRITE_BACK IS
	GENERIC (
		CELL_SIZE : INTEGER := 4;
		MEMORY_ADDRESS_WIDTH : INTEGER := 27;
		NUMBER_OF_ROWS : INTEGER := 1080; -- FOR EXAMPLE: 1080 FOR 1080 LINES
		NEIGHBORHOOD_SIZE : INTEGER := 5; -- FOR EXAMPLE: 7 FOR AN 7X7 NEIGHBORHOOD
		GRID_TYPE : STRING  := "TOROIDAL"; 
		-- VALID VALUES: "RECTANGULAR", "CYLINDRICAL" AND "TOROIDAL"
		NUMBER_OF_BURSTS_PER_LINE : INTEGER := 60; -- 
		BURST_SIZE : INTEGER := 128;
		SPEED : INTEGER := 120
	);
	PORT ( 	
		CLK : IN STD_LOGIC;	-- UI_CLK FROM MIG DDR CONTROLLER
		RST : IN STD_LOGIC;
		-- CONTROL SIGNALS --
		MEM_ACCESS_GRANTED : IN STD_LOGIC;
		-- FIFO SIGNALS
		FIFO_DATA : IN STD_LOGIC_VECTOR(BURST_SIZE-1 DOWNTO 0);
		FIFO_READ_EN : OUT STD_LOGIC := '0';
		FIFO_READY : IN STD_LOGIC; -- FIFO_READY = NOT EMPTY
		-- 
		SPEED_SETTING : IN INTEGER RANGE 0 TO SPEED; -- GRAPHICS RUN AT 60 FPS. SPEED = 60: NEW GENERATION EVERY 1 SEC. SPEED = 0: FULL SPEED, NEW GENERATION EVERY NEW FRAME.
		WB_SPEED_COUNTER : OUT INTEGER RANGE 0 TO SPEED := 0;
		--
		COLUMN_BEING_WRITTEN : OUT INTEGER RANGE 0 TO NUMBER_OF_BURSTS_PER_LINE;
		ROW_BEING_WRITTEN : OUT INTEGER RANGE 0 TO NUMBER_OF_ROWS-1;
		-- MEMORY SIGNALS --
		APP_RDY : IN STD_LOGIC;
		APP_WDF_RDY : IN STD_LOGIC;
		APP_EN : OUT STD_LOGIC := '0';
		APP_CMD : OUT STD_LOGIC_VECTOR(2 DOWNTO 0) := "000"; -- "000" = WRITE COMMAND
		APP_WDF_DATA : OUT STD_LOGIC_VECTOR(BURST_SIZE-1 DOWNTO 0);
		APP_WDF_END : OUT STD_LOGIC := '0';
		APP_WDF_WREN : OUT STD_LOGIC := '0';
		APP_ADDR : OUT STD_LOGIC_VECTOR(MEMORY_ADDRESS_WIDTH-1 DOWNTO 0)
	);
END WRITE_BACK;

ARCHITECTURE BEHAVIORAL OF WRITE_BACK IS	
	
	-- TOROIDAL GRID: GRID_X x GRID_Y cells
	-- RECT OR CYLINDR GRID: GRID_X x (GRID_Y-(NEIGHBORHOOD_SIZE-1)) cells
	function init return INTEGER is
	begin
		IF (GRID_TYPE = "TOROIDAL") THEN
			return 0;
		ELSE
			return (NEIGHBORHOOD_SIZE-1)/2;
		END IF;
	end function init;
	
	SIGNAL ADDRESS_COLUMN : INTEGER RANGE 0 TO NUMBER_OF_BURSTS_PER_LINE := 0;
	SIGNAL BURSTS_RECEIVED_FROM_FIFO_COUNTER, BURSTS_WRITTEN_COUNTER, COMMANDS_SENT_COUNTER : INTEGER RANGE 0 TO NUMBER_OF_BURSTS_PER_LINE := 0;
	SIGNAL ADDRESS_ROW : INTEGER RANGE 0 TO NUMBER_OF_ROWS-1 := init;
	SIGNAL SPEED_COUNTER : INTEGER RANGE 0 TO SPEED := 0;
	SIGNAL APP_WDF_WREN_SIGNAL, APP_WDF_END_SIGNAL, APP_EN_SIGNAL : STD_LOGIC := '0';
	
	SIGNAL SELECTED_FRAME : STD_LOGIC := '1';
	
	constant ADDRESS_ROW_INIT : INTEGER := init;
	
BEGIN

	-- THE FOLLOWING FSM HANDLES THE DATA BEING RECEIVED  
	WRITE_MEMORY: PROCESS 
	BEGIN
		
		WAIT UNTIL RISING_EDGE(CLK);
		
		IF RST = '1' THEN
			ADDRESS_COLUMN <= 0;
			ADDRESS_ROW <= ADDRESS_ROW_INIT;
			APP_WDF_WREN_SIGNAL <= '0';
			APP_WDF_END_SIGNAL <= '0';
			SELECTED_FRAME <= '1';
			BURSTS_RECEIVED_FROM_FIFO_COUNTER <= 0;
			BURSTS_WRITTEN_COUNTER <= 0;
			COMMANDS_SENT_COUNTER <= 0;
			SPEED_COUNTER <= 0;
		ELSE
			IF APP_EN_SIGNAL = '1' AND APP_RDY = '1' THEN
				IF ADDRESS_COLUMN = NUMBER_OF_BURSTS_PER_LINE-1 THEN
					ADDRESS_COLUMN <= 0;
					-- CHANGE LINE
					IF ADDRESS_ROW = (NUMBER_OF_ROWS-1)-ADDRESS_ROW_INIT THEN 
						IF SPEED_COUNTER >= SPEED_SETTING THEN
							SPEED_COUNTER <= 0;
							SELECTED_FRAME <= NOT SELECTED_FRAME;
						ELSE
							IF SPEED_SETTING = SPEED-1 THEN -- SIM ENDED
								 SPEED_COUNTER <= SPEED_COUNTER;
							ELSE	 
								 SPEED_COUNTER <= SPEED_COUNTER + 1;
							END IF;
						END IF;
						ADDRESS_ROW <= ADDRESS_ROW_INIT;
					ELSE	
						ADDRESS_ROW <= ADDRESS_ROW + 1;
					END IF;
				ELSE
					ADDRESS_COLUMN <= ADDRESS_COLUMN + 1;
				END IF;
				
				IF COMMANDS_SENT_COUNTER = NUMBER_OF_BURSTS_PER_LINE-1 THEN
					COMMANDS_SENT_COUNTER <= 0;
					BURSTS_WRITTEN_COUNTER <= 0;
					BURSTS_RECEIVED_FROM_FIFO_COUNTER <= 0;
				ELSE
					COMMANDS_SENT_COUNTER <= COMMANDS_SENT_COUNTER + 1;
				END IF;
				
			END IF;
			
			-- IF BURSTS_WRITTEN_COUNTER > COMMANDS_SENT_COUNTER AND APP_RDY = '1' THEN
				-- APP_EN_SIGNAL <= '1';
			-- ELSE
				-- APP_EN_SIGNAL <= '0';
			-- END IF;
			
			IF APP_WDF_RDY = '1' AND (APP_WDF_WREN_SIGNAL = '1' OR (BURSTS_RECEIVED_FROM_FIFO_COUNTER > BURSTS_WRITTEN_COUNTER AND APP_WDF_RDY = '1')) AND MEM_ACCESS_GRANTED = '1' THEN 
				BURSTS_WRITTEN_COUNTER <= BURSTS_WRITTEN_COUNTER + 1;
			END IF;
			
			IF FIFO_READY = '1' AND APP_WDF_RDY = '1' AND MEM_ACCESS_GRANTED = '1' THEN
				APP_WDF_WREN_SIGNAL <= '1';
				APP_WDF_END_SIGNAL <= '1';
				--------------------------------------------------------------------------
				BURSTS_RECEIVED_FROM_FIFO_COUNTER <= BURSTS_RECEIVED_FROM_FIFO_COUNTER + 1;
				--------------------------------------------------------------------------
			ELSE
				APP_WDF_WREN_SIGNAL <= '0';
				APP_WDF_END_SIGNAL <= '0';
			END IF;
		END IF;
	END PROCESS WRITE_MEMORY;
	
	PROCESS(FIFO_DATA)
	BEGIN
		-- NOT TO BE CONFUSED WITH 
		-- APP_WDF_DATA( ((31-i+1)*CELL_SIZE)-1 DOWNTO (31 - i)*CELL_SIZE )
		IF CELL_SIZE = 4 THEN
			for i in 0 to 31 loop
				APP_WDF_DATA( ((31-i+1)*4)-1 DOWNTO (31 - i)*4 ) <= FIFO_DATA ( ((i+1)*4)-1 DOWNTO i*4 );
			end loop ; 
		ELSE
			for i in 0 to 15 loop
				APP_WDF_DATA( ((15-i+1)*8)-1 DOWNTO (15 - i)*8 ) <= FIFO_DATA ( ((i+1)*8)-1 DOWNTO i*8 ) ;
			end loop;
		END IF; 
	END PROCESS;
	
	FIFO_READ_EN <= APP_WDF_RDY WHEN FIFO_READY = '1' AND MEM_ACCESS_GRANTED = '1' ELSE '0';
	
	APP_EN_SIGNAL <= '1' WHEN BURSTS_WRITTEN_COUNTER > COMMANDS_SENT_COUNTER AND APP_RDY = '1' ELSE '0';
	APP_EN <= '1' WHEN BURSTS_WRITTEN_COUNTER > COMMANDS_SENT_COUNTER AND APP_RDY = '1' ELSE '0'; -- APP EN SIGNAL
	
	-- APP_WDF_WREN <= APP_WDF_WREN_SIGNAL;
	-- APP_WDF_END <= APP_WDF_END_SIGNAL;
	APP_WDF_WREN <= '1' WHEN APP_WDF_WREN_SIGNAL = '1' OR (BURSTS_RECEIVED_FROM_FIFO_COUNTER > BURSTS_WRITTEN_COUNTER AND APP_WDF_RDY = '1') ELSE '0';
	APP_WDF_END <= '1' WHEN APP_WDF_END_SIGNAL = '1' OR (BURSTS_RECEIVED_FROM_FIFO_COUNTER > BURSTS_WRITTEN_COUNTER AND APP_WDF_RDY = '1') ELSE '0';
	
	APP_ADDR(19 DOWNTO 0) <= STD_LOGIC_VECTOR(TO_UNSIGNED((ADDRESS_ROW*NUMBER_OF_BURSTS_PER_LINE*8 ) + ADDRESS_COLUMN*8, 20));
	APP_ADDR(20) <= SELECTED_FRAME;
	APP_ADDR(MEMORY_ADDRESS_WIDTH-1 DOWNTO 21) <= (OTHERS => '0');
	
	COLUMN_BEING_WRITTEN <= BURSTS_WRITTEN_COUNTER;
	ROW_BEING_WRITTEN <= ADDRESS_ROW;

	APP_CMD <= "000"; -- WRITE COMMAND
	
	WB_SPEED_COUNTER <= SPEED_COUNTER;

END BEHAVIORAL;